`include "fifomemory.v"
module fifomemory_tb;
parameter DEPTH=16;
parameter PTR_WIDTH=$clog2(DEPTH);
parameter WIDTH=8;
reg clk_i,rst_i;
reg wr_en_i,rd_en_i;
reg [WIDTH-1:0]wdata_i;
wire [WIDTH-1:0]rdata_o;
wire wr_error_o,rd_error_o;
wire full_o,empty_o;
reg [WIDTH-1:0]mem[DEPTH-1:0];
//reg [PTR_WIDTH-1:0]wr_ptr;
//reg [PTR_WIDTH-1:0]rd_ptr;
//reg wr_toggle_f,rd_toggle_f;
integer i;
fifomemory dut(clk_i,rst_i,wr_en_i,wdata_i,rd_en_i,rdata_o,full_o,empty_o,wr_error_o,rd_error_o);
initial begin
	clk_i=0;
	forever #5 clk_i=~clk_i;
end
initial begin
	reset_fifo();
	write_fifo(DEPTH);
	read_fifo(DEPTH);
end	
task reset_fifo();
begin
	rst_i=1;
	wr_en_i=0;
	rd_en_i=0;
	wdata_i=0;
	@(posedge clk_i);
	rst_i=0;
end
endtask
task write_fifo(input integer num_loc);
begin
	for(i=0;i<num_loc;i=i+1)begin
		@(posedge clk_i);
		wr_en_i=1;
		wdata_i=$random;
	end
		@(posedge clk_i);
		wr_en_i=0;
		wdata_i=0;
end
endtask
task read_fifo(input integer num_loc);
begin
	for(i=0;i<num_loc;i=i+1)begin
		@(posedge clk_i);
			rd_en_i=1;
	end
		@(posedge clk_i);
			rd_en_i=0;
end
endtask
initial begin
	#1000;
	$finish;
end	
endmodule
