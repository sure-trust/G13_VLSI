module ha(a,b,s,c);
input a,b;
input s,c;
assign s=a^b;
assign c=a&b;
endmodule 


